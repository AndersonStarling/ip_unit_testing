`timescale 1ns / 1ps



module test_flip_flop();





endmodule